module uart(
);
endmodule